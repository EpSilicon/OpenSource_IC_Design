magic
tech sky130A
magscale 1 2
timestamp 1711820162
<< nmos >>
rect -229 -4000 -29 4000
rect 29 -4000 229 4000
<< ndiff >>
rect -287 3988 -229 4000
rect -287 -3988 -275 3988
rect -241 -3988 -229 3988
rect -287 -4000 -229 -3988
rect -29 3988 29 4000
rect -29 -3988 -17 3988
rect 17 -3988 29 3988
rect -29 -4000 29 -3988
rect 229 3988 287 4000
rect 229 -3988 241 3988
rect 275 -3988 287 3988
rect 229 -4000 287 -3988
<< ndiffc >>
rect -275 -3988 -241 3988
rect -17 -3988 17 3988
rect 241 -3988 275 3988
<< poly >>
rect -229 4072 -29 4088
rect -229 4038 -213 4072
rect -45 4038 -29 4072
rect -229 4000 -29 4038
rect 29 4072 229 4088
rect 29 4038 45 4072
rect 213 4038 229 4072
rect 29 4000 229 4038
rect -229 -4038 -29 -4000
rect -229 -4072 -213 -4038
rect -45 -4072 -29 -4038
rect -229 -4088 -29 -4072
rect 29 -4038 229 -4000
rect 29 -4072 45 -4038
rect 213 -4072 229 -4038
rect 29 -4088 229 -4072
<< polycont >>
rect -213 4038 -45 4072
rect 45 4038 213 4072
rect -213 -4072 -45 -4038
rect 45 -4072 213 -4038
<< locali >>
rect -229 4038 -213 4072
rect -45 4038 -29 4072
rect 29 4038 45 4072
rect 213 4038 229 4072
rect -275 3988 -241 4004
rect -275 -4004 -241 -3988
rect -17 3988 17 4004
rect -17 -4004 17 -3988
rect 241 3988 275 4004
rect 241 -4004 275 -3988
rect -229 -4072 -213 -4038
rect -45 -4072 -29 -4038
rect 29 -4072 45 -4038
rect 213 -4072 229 -4038
<< viali >>
rect -213 4038 -45 4072
rect 45 4038 213 4072
rect -275 -3988 -241 3988
rect -17 -3988 17 3988
rect 241 -3988 275 3988
rect -213 -4072 -45 -4038
rect 45 -4072 213 -4038
<< metal1 >>
rect -225 4072 -33 4078
rect -225 4038 -213 4072
rect -45 4038 -33 4072
rect -225 4032 -33 4038
rect 33 4072 225 4078
rect 33 4038 45 4072
rect 213 4038 225 4072
rect 33 4032 225 4038
rect -281 3988 -235 4000
rect -281 -3988 -275 3988
rect -241 -3988 -235 3988
rect -281 -4000 -235 -3988
rect -23 3988 23 4000
rect -23 -3988 -17 3988
rect 17 -3988 23 3988
rect -23 -4000 23 -3988
rect 235 3988 281 4000
rect 235 -3988 241 3988
rect 275 -3988 281 3988
rect 235 -4000 281 -3988
rect -225 -4038 -33 -4032
rect -225 -4072 -213 -4038
rect -45 -4072 -33 -4038
rect -225 -4078 -33 -4072
rect 33 -4038 225 -4032
rect 33 -4072 45 -4038
rect 213 -4072 225 -4038
rect 33 -4078 225 -4072
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 40.0 l 1.0 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
