magic
tech sky130A
magscale 1 2
timestamp 1711887509
<< locali >>
rect 10247 7063 10364 7098
rect 10254 6677 10371 6712
rect 10247 6291 10364 6325
rect 12338 4688 12462 4722
rect 12338 4202 12462 4236
rect 12338 3716 12462 3750
rect 12338 3230 12462 3264
<< viali >>
rect 6172 7335 10345 7369
rect 4272 3116 12366 3150
<< metal1 >>
rect 4117 7369 10371 7504
rect 4117 7335 6172 7369
rect 10345 7335 10371 7369
rect 4117 7297 10371 7335
rect 6172 7215 6271 7261
rect 8336 7258 8460 7268
rect 6172 7193 6218 7215
rect 8336 7206 8346 7258
rect 8450 7206 8460 7258
rect 8336 7196 8460 7206
rect 6177 6726 6211 7193
rect 8940 6884 9064 6892
rect 8940 6832 8948 6884
rect 9052 6832 9064 6884
rect 8940 6828 9064 6832
rect 6258 6634 12585 6643
rect 6258 6504 9570 6634
rect 9666 6504 12585 6634
rect 6258 6443 12585 6504
rect 6177 6342 6211 6432
rect 6170 6332 9060 6342
rect 6170 6266 8952 6332
rect 9048 6266 9060 6332
rect 6170 6258 9060 6266
rect 8334 5970 8460 5980
rect 8334 5918 8346 5970
rect 8448 5918 8460 5970
rect 8334 5906 8460 5918
rect 4120 5706 4320 5906
rect 7726 5696 7846 5706
rect 7726 5644 7736 5696
rect 7838 5644 7846 5696
rect 7726 5636 7846 5644
rect 8942 5480 9062 5486
rect 8942 5428 8948 5480
rect 9056 5428 9062 5480
rect 8942 5426 9062 5428
rect 4120 5220 4320 5420
rect 7724 5210 7848 5218
rect 7724 5158 7736 5210
rect 7838 5158 7848 5210
rect 7724 5150 7848 5158
rect 7726 4996 7846 5004
rect 7726 4944 7734 4996
rect 7838 4944 7846 4996
rect 7726 4934 7846 4944
rect 4272 3528 4320 4930
rect 7724 4508 7850 4516
rect 7724 4456 7732 4508
rect 7842 4456 7850 4508
rect 7724 4448 7850 4456
rect 9558 4022 9680 4028
rect 9558 3970 9564 4022
rect 9674 3970 9680 4022
rect 9558 3968 9680 3970
rect 4272 3482 4454 3528
rect 4272 3476 4320 3482
rect 4120 3276 4320 3476
rect 4120 3150 12466 3160
rect 4120 3116 4272 3150
rect 12366 3116 12466 3150
rect 4120 2960 12466 3116
<< via1 >>
rect 8346 7206 8450 7258
rect 8948 6832 9052 6884
rect 9570 6504 9666 6634
rect 8952 6266 9048 6332
rect 8346 5918 8448 5970
rect 7736 5644 7838 5696
rect 8948 5428 9056 5480
rect 7736 5158 7838 5210
rect 7734 4944 7838 4996
rect 7732 4456 7842 4508
rect 9564 3970 9674 4022
<< metal2 >>
rect 8336 7258 8460 7268
rect 8336 7206 8346 7258
rect 8450 7206 8460 7258
rect 8336 7196 8460 7206
rect 8341 5980 8455 7196
rect 8945 6884 9059 6892
rect 8945 6832 8948 6884
rect 9052 6832 9059 6884
rect 8945 6332 9059 6832
rect 8945 6266 8952 6332
rect 9048 6266 9059 6332
rect 8334 5970 8460 5980
rect 8334 5918 8346 5970
rect 8448 5918 8460 5970
rect 8334 5906 8460 5918
rect 7726 5696 7846 5706
rect 7726 5644 7736 5696
rect 7838 5644 7846 5696
rect 7726 5636 7846 5644
rect 7730 5218 7844 5636
rect 8945 5480 9059 6266
rect 8945 5428 8948 5480
rect 9056 5428 9059 5480
rect 8945 5420 9059 5428
rect 9563 6634 9677 6642
rect 9563 6504 9570 6634
rect 9666 6504 9677 6634
rect 7724 5210 7848 5218
rect 7724 5158 7736 5210
rect 7838 5158 7848 5210
rect 7724 5150 7848 5158
rect 7730 5004 7844 5150
rect 7726 4996 7846 5004
rect 7726 4944 7734 4996
rect 7838 4944 7846 4996
rect 7726 4934 7846 4944
rect 7730 4516 7844 4934
rect 7724 4508 7850 4516
rect 7724 4456 7732 4508
rect 7842 4456 7850 4508
rect 7724 4448 7850 4456
rect 9563 4022 9677 6504
rect 9563 3970 9564 4022
rect 9674 3970 9677 4022
rect 9563 3962 9677 3970
use sky130_fd_pr__nfet_01v8  sky130_fd_pr__nfet_01v8_0
timestamp 1711887509
transform 1 0 2236 0 1 -3060
box 0 0 1 1
use sky130_fd_pr__nfet_01v8  sky130_fd_pr__nfet_01v8_1
timestamp 1711887509
transform 1 0 2237 0 1 -3060
box 0 0 1 1
use sky130_fd_pr__nfet_01v8_KWM3S5  sky130_fd_pr__nfet_01v8_KWM3S5_0
timestamp 1711879029
transform 0 1 8319 -1 0 3376
box -296 -4179 296 4179
use sky130_fd_pr__pfet_01v8_LZG3QU  sky130_fd_pr__pfet_01v8_LZG3QU_0
timestamp 1711879029
transform 0 1 8223 -1 0 6773
box -246 -2184 246 2184
use sky130_fd_pr__pfet_01v8_LZG3QU  sky130_fd_pr__pfet_01v8_LZG3QU_1
timestamp 1711879029
transform 0 1 8223 -1 0 6387
box -246 -2184 246 2184
use sky130_fd_pr__nfet_01v8_K2PRWZ  XM1
timestamp 1711879029
transform 0 1 8319 -1 0 5806
box -296 -4179 296 4179
use sky130_fd_pr__nfet_01v8_K2PRWZ  XM2
timestamp 1711879029
transform 0 1 8319 -1 0 5320
box -296 -4179 296 4179
use sky130_fd_pr__pfet_01v8_LZG3QU  XM3
timestamp 1711879029
transform 0 1 8223 -1 0 7159
box -246 -2184 246 2184
use sky130_fd_pr__nfet_01v8  XM6[0]
timestamp 1711887509
transform 1 0 2396 0 1 -3325
box 0 0 1 1
use sky130_fd_pr__nfet_01v8  XM6[1]
timestamp 1711887509
transform 1 0 2395 0 1 -3325
box 0 0 1 1
use sky130_fd_pr__nfet_01v8_KWM3S5  XM6_0
timestamp 1711879029
transform 0 1 8319 -1 0 4348
box -296 -4179 296 4179
use sky130_fd_pr__nfet_01v8_KWM3S5  XM6_1
timestamp 1711879029
transform 0 1 8319 -1 0 4834
box -296 -4179 296 4179
use sky130_fd_pr__nfet_01v8_KWM3S5  XM7
timestamp 1711879029
transform 0 1 8319 -1 0 3862
box -296 -4179 296 4179
<< labels >>
flabel metal1 4120 5706 4320 5906 0 FreeSans 256 0 0 0 inn
port 3 nsew
flabel metal1 4120 5220 4320 5420 0 FreeSans 256 0 0 0 inp
port 2 nsew
flabel metal1 4120 3276 4320 3476 0 FreeSans 256 0 0 0 ibiasn
port 4 nsew
flabel metal1 4120 7300 4320 7500 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 12385 6443 12585 6643 0 FreeSans 256 0 0 0 out
port 1 nsew
flabel metal1 4120 2960 4320 3160 0 FreeSans 256 0 0 0 vss
port 5 nsew
<< end >>
