* NGSPICE file created from opamp.ext - technology: sky130A

.subckt opamp_ext_RC vdd out inp inn ibiasn vss
X0 vss ibiasn ibiasn vss sky130_fd_pr__nfet_01v8 ad=11.6 pd=80.58 as=11.6 ps=80.58 w=40 l=1
X1 m1_7724_4448# inn m1_8334_5906# vss sky130_fd_pr__nfet_01v8 ad=11.6 pd=80.58 as=11.6 ps=80.58 w=40 l=1
X2 m1_7724_4448# inp m1_6170_6258# vss sky130_fd_pr__nfet_01v8 ad=11.6 pd=80.58 as=11.6 ps=80.58 w=40 l=1
X3 vdd m1_8334_5906# m1_8334_5906# vdd sky130_fd_pr__pfet_01v8 ad=5.8 pd=40.58 as=5.8 ps=40.58 w=20 l=0.5
X4 vss ibiasn m1_7724_4448# vss sky130_fd_pr__nfet_01v8 ad=11.6 pd=80.58 as=11.6 ps=80.58 w=40 l=1
X5 vss ibiasn m1_7724_4448# vss sky130_fd_pr__nfet_01v8 ad=11.6 pd=80.58 as=11.6 ps=80.58 w=40 l=1
X6 vss ibiasn out vss sky130_fd_pr__nfet_01v8 ad=11.6 pd=80.58 as=11.6 ps=80.58 w=40 l=1
X7 vdd m1_8334_5906# m1_6170_6258# vdd sky130_fd_pr__pfet_01v8 ad=5.8 pd=40.58 as=5.8 ps=40.58 w=20 l=0.5
X8 vdd m1_6170_6258# out vdd sky130_fd_pr__pfet_01v8 ad=5.8 pd=40.58 as=5.8 ps=40.58 w=20 l=0.5
C0 inp m1_8334_5906# 0.002675f
C1 inn m1_7724_4448# 0.867763f
C2 ibiasn m1_6170_6258# 0.003701f
C3 out inn 0.07251f
C4 m1_8334_5906# m1_7724_4448# 2.189434f
C5 vdd m1_6170_6258# 3.070694f
C6 m1_8334_5906# out 0.818384f
C7 inp m1_7724_4448# 0.944646f
C8 inp out 0.083426f
C9 inn m1_6170_6258# 0.072016f
C10 out m1_7724_4448# 1.118943f
C11 m1_8334_5906# m1_6170_6258# 1.717438f
C12 inp m1_6170_6258# 0.867091f
C13 m1_6170_6258# m1_7724_4448# 3.938311f
C14 vdd inn 0.00629f
C15 ibiasn m1_8334_5906# 0.001415f
C16 out m1_6170_6258# 2.295279f
C17 m1_8334_5906# vdd 4.940537f
C18 ibiasn inp 0.013092f
C19 ibiasn m1_7724_4448# 2.187538f
C20 ibiasn out 2.139875f
C21 m1_8334_5906# inn 0.868036f
C22 vdd m1_7724_4448# 0.003134f
C23 vdd out 2.937594f
C24 inp inn 0.032568f
R0 ibiasn.n0 ibiasn.t3 1059.17
R1 ibiasn.n3 ibiasn.t0 1057.91
R2 ibiasn.n0 ibiasn.t2 1057.91
R3 ibiasn.n1 ibiasn.t4 1057.91
R4 ibiasn.n2 ibiasn.t1 13.0516
R5 ibiasn.n1 ibiasn.n0 1.26612
R6 ibiasn.n2 ibiasn.n1 0.930188
R7 ibiasn.n3 ibiasn.n2 0.138521
R8 ibiasn ibiasn.n3 0.063
R9 vss.n59 vss.n1 25216
R10 vss.n38 vss.n1 25216
R11 vss.n31 vss.n9 25216
R12 vss.n57 vss.n9 25216
R13 vss.n37 vss.n17 23906.5
R14 vss.n17 vss.n3 23906.5
R15 vss.n49 vss.n21 23906.5
R16 vss.n49 vss.n22 23906.5
R17 vss.n25 vss.n19 23906.5
R18 vss.n19 vss.n18 23906.5
R19 vss.n51 vss.n15 23906.5
R20 vss.n51 vss.n16 23906.5
R21 vss.n32 vss.n20 23906.5
R22 vss.n20 vss.n10 23906.5
R23 vss.n39 vss.n4 5520.18
R24 vss.n58 vss.n4 5516.42
R25 vss.n56 vss.n11 1638.4
R26 vss.n33 vss.n11 1638.4
R27 vss.n61 vss.n60 1638.4
R28 vss.n61 vss.n0 1625.6
R29 vss.n34 vss.n12 1553.32
R30 vss.n55 vss.n12 1553.32
R31 vss.n52 vss.n14 1553.32
R32 vss.n53 vss.n52 1553.32
R33 vss.n43 vss.n42 1553.32
R34 vss.n44 vss.n43 1553.32
R35 vss.n48 vss.n23 1553.32
R36 vss.n48 vss.n47 1553.32
R37 vss.n27 vss.n26 1553.32
R38 vss.n26 vss.n2 1553.32
R39 vss.n59 vss.n3 1309.47
R40 vss.n29 vss.n21 1309.47
R41 vss.n37 vss.n29 1309.47
R42 vss.n38 vss.n37 1309.47
R43 vss.n18 vss.n6 1309.47
R44 vss.n22 vss.n6 1309.47
R45 vss.n22 vss.n5 1309.47
R46 vss.n5 vss.n3 1309.47
R47 vss.n30 vss.n15 1309.47
R48 vss.n30 vss.n25 1309.47
R49 vss.n40 vss.n25 1309.47
R50 vss.n40 vss.n21 1309.47
R51 vss.n10 vss.n8 1309.47
R52 vss.n16 vss.n8 1309.47
R53 vss.n16 vss.n7 1309.47
R54 vss.n18 vss.n7 1309.47
R55 vss.n32 vss.n31 1309.47
R56 vss.n36 vss.n32 1309.47
R57 vss.n36 vss.n15 1309.47
R58 vss.n57 vss.n10 1309.47
R59 vss.n57 vss.n56 117.001
R60 vss.n58 vss.n57 117.001
R61 vss.n33 vss.n31 117.001
R62 vss.n39 vss.n31 117.001
R63 vss.n36 vss.n35 117.001
R64 vss.n39 vss.n36 117.001
R65 vss.n54 vss.n8 117.001
R66 vss.n58 vss.n8 117.001
R67 vss.n13 vss.n7 117.001
R68 vss.n58 vss.n7 117.001
R69 vss.n30 vss.n24 117.001
R70 vss.n39 vss.n30 117.001
R71 vss.n41 vss.n40 117.001
R72 vss.n40 vss.n39 117.001
R73 vss.n45 vss.n6 117.001
R74 vss.n58 vss.n6 117.001
R75 vss.n46 vss.n5 117.001
R76 vss.n58 vss.n5 117.001
R77 vss.n29 vss.n28 117.001
R78 vss.n39 vss.n29 117.001
R79 vss.n38 vss.n0 117.001
R80 vss.n39 vss.n38 117.001
R81 vss.n60 vss.n59 117.001
R82 vss.n59 vss.n58 117.001
R83 vss.n50 vss.n4 94.4106
R84 vss.n56 vss.n55 85.0829
R85 vss.n34 vss.n33 85.0829
R86 vss.n35 vss.n34 85.0829
R87 vss.n35 vss.n14 85.0829
R88 vss.n55 vss.n54 85.0829
R89 vss.n54 vss.n53 85.0829
R90 vss.n53 vss.n13 85.0829
R91 vss.n44 vss.n13 85.0829
R92 vss.n24 vss.n14 85.0829
R93 vss.n42 vss.n41 85.0829
R94 vss.n45 vss.n44 85.0829
R95 vss.n47 vss.n45 85.0829
R96 vss.n47 vss.n46 85.0829
R97 vss.n46 vss.n2 85.0829
R98 vss.n28 vss.n23 85.0829
R99 vss.n27 vss.n0 85.0829
R100 vss.n60 vss.n2 85.0829
R101 vss.n41 vss.n23 72.2828
R102 vss.n42 vss.n24 72.2828
R103 vss.n28 vss.n27 72.2828
R104 vss.n11 vss.n9 4.91647
R105 vss.n50 vss.n9 4.91647
R106 vss.n20 vss.n12 4.91647
R107 vss.n50 vss.n20 4.91647
R108 vss.n52 vss.n51 4.91647
R109 vss.n51 vss.n50 4.91647
R110 vss.n43 vss.n19 4.91647
R111 vss.n50 vss.n19 4.91647
R112 vss.n49 vss.n48 4.91647
R113 vss.n50 vss.n49 4.91647
R114 vss.n26 vss.n17 4.91647
R115 vss.n50 vss.n17 4.91647
R116 vss.n61 vss.n1 4.91647
R117 vss.n50 vss.n1 4.91647
R118 vss vss.n61 2.70791
R119 inn inn.t0 1058.01
R120 inp inp.t0 1058.01
R121 vdd.n20 vdd.n6 8142.35
R122 vdd.n23 vdd.n6 8142.35
R123 vdd.n29 vdd.n2 8142.35
R124 vdd.n29 vdd.n3 8142.35
R125 vdd.n27 vdd.n8 7521.18
R126 vdd.n27 vdd.n9 7521.18
R127 vdd.n11 vdd.n5 7521.18
R128 vdd.n17 vdd.n5 7521.18
R129 vdd.n28 vdd.n4 1601.62
R130 vdd.n28 vdd.n7 1601.62
R131 vdd.n24 vdd.n22 868.519
R132 vdd.n30 vdd.n1 868.519
R133 vdd.n22 vdd.n21 855.718
R134 vdd.n31 vdd.n0 855.341
R135 vdd.n26 vdd.n10 802.26
R136 vdd.n26 vdd.n25 802.26
R137 vdd.n15 vdd.n14 802.26
R138 vdd.n16 vdd.n15 802.26
R139 vdd.n20 vdd.n8 621.178
R140 vdd.n18 vdd.n17 621.178
R141 vdd.n18 vdd.n9 621.178
R142 vdd.n23 vdd.n9 621.178
R143 vdd.n11 vdd.n2 621.178
R144 vdd.n12 vdd.n11 621.178
R145 vdd.n12 vdd.n8 621.178
R146 vdd.n17 vdd.n3 621.178
R147 vdd.n14 vdd.n13 66.2593
R148 vdd.n25 vdd.n24 66.2593
R149 vdd.n21 vdd.n10 66.2593
R150 vdd.n16 vdd.n1 66.2593
R151 vdd.n19 vdd.n16 66.2593
R152 vdd.n25 vdd.n19 66.2593
R153 vdd.n21 vdd.n20 61.6672
R154 vdd.n20 vdd.n4 61.6672
R155 vdd.n24 vdd.n23 61.6672
R156 vdd.n23 vdd.n7 61.6672
R157 vdd.n13 vdd.n12 61.6672
R158 vdd.n12 vdd.n4 61.6672
R159 vdd.n3 vdd.n1 61.6672
R160 vdd.n7 vdd.n3 61.6672
R161 vdd.n19 vdd.n18 61.6672
R162 vdd.n18 vdd.n7 61.6672
R163 vdd.n2 vdd.n0 61.6672
R164 vdd.n4 vdd.n2 61.6672
R165 vdd.n13 vdd.n10 53.0829
R166 vdd.n14 vdd.n0 53.0829
R167 vdd.n31 vdd.n30 13.177
R168 vdd.n22 vdd.n6 3.08383
R169 vdd.n28 vdd.n6 3.08383
R170 vdd.n27 vdd.n26 3.08383
R171 vdd.n28 vdd.n27 3.08383
R172 vdd.n15 vdd.n5 3.08383
R173 vdd.n28 vdd.n5 3.08383
R174 vdd.n30 vdd.n29 3.08383
R175 vdd.n29 vdd.n28 3.08383
R176 vdd vdd.n31 2.65964
C25 vdd.n1 vss 0.059365f
C26 vdd.n2 vss 0.059365f
C27 vdd.n3 vss 0.059365f
C28 vdd.n4 vss 1.96349f
C29 vdd.n5 vss 0.100626f
C30 vdd.n6 vss 0.109059f
C31 vdd.n7 vss 1.96349f
C32 vdd.n8 vss 0.059426f
C33 vdd.n9 vss 0.059426f
C34 vdd.n10 vss 0.00336f
C35 vdd.n11 vss 0.059426f
C36 vdd.n12 vss 0.008311f
C37 vdd.n14 vss 0.003363f
C38 vdd.n15 vss 0.100626f
C39 vdd.n16 vss 0.059426f
C40 vdd.n17 vss 0.059426f
C41 vdd.n18 vss 0.008311f
C42 vdd.n19 vss 0.008311f
C43 vdd.n20 vss 0.059365f
C44 vdd.n22 vss 0.104758f
C45 vdd.n23 vss 0.059365f
C46 vdd.n24 vss 0.059365f
C47 vdd.n25 vss 0.059426f
C48 vdd.n26 vss 0.100626f
C49 vdd.n27 vss 0.100626f
C50 vdd.n28 vss 3.7409f
C51 vdd.n29 vss 0.109059f
C52 vdd.n30 vss 0.055356f
C53 vdd.n31 vss 1.1843f
C54 ibiasn.t1 vss 0.511366f
C55 ibiasn.t3 vss 0.688822f
C56 ibiasn.t2 vss 0.688552f
C57 ibiasn.n0 vss 0.455043f
C58 ibiasn.t4 vss 0.688552f
C59 ibiasn.n1 vss 0.227898f
C60 ibiasn.n2 vss 0.114584f
C61 ibiasn.t0 vss 0.688552f
C62 ibiasn.n3 vss 0.23104f
C63 out vss 14.865181f
C64 ibiasn vss 10.046253f
C65 m1_7724_4448# vss 20.980135f
C66 m1_8334_5906# vss 5.273708f
C67 vdd vss 23.929913f
C68 m1_6170_6258# vss 5.563833f
C69 inp vss 0.601188f
C70 inn vss 0.606819f
.ends
