magic
tech sky130A
timestamp 1711887509
<< end >>
