magic
tech sky130A
magscale 1 2
timestamp 1711820162
<< nwell >>
rect -325 -2219 325 2219
<< pmos >>
rect -129 -2000 -29 2000
rect 29 -2000 129 2000
<< pdiff >>
rect -187 1988 -129 2000
rect -187 -1988 -175 1988
rect -141 -1988 -129 1988
rect -187 -2000 -129 -1988
rect -29 1988 29 2000
rect -29 -1988 -17 1988
rect 17 -1988 29 1988
rect -29 -2000 29 -1988
rect 129 1988 187 2000
rect 129 -1988 141 1988
rect 175 -1988 187 1988
rect 129 -2000 187 -1988
<< pdiffc >>
rect -175 -1988 -141 1988
rect -17 -1988 17 1988
rect 141 -1988 175 1988
<< nsubdiff >>
rect -289 2149 -193 2183
rect 193 2149 289 2183
rect -289 2087 -255 2149
rect 255 2087 289 2149
rect -289 -2149 -255 -2087
rect 255 -2149 289 -2087
rect -289 -2183 -193 -2149
rect 193 -2183 289 -2149
<< nsubdiffcont >>
rect -193 2149 193 2183
rect -289 -2087 -255 2087
rect 255 -2087 289 2087
rect -193 -2183 193 -2149
<< poly >>
rect -129 2081 -29 2097
rect -129 2047 -113 2081
rect -45 2047 -29 2081
rect -129 2000 -29 2047
rect 29 2081 129 2097
rect 29 2047 45 2081
rect 113 2047 129 2081
rect 29 2000 129 2047
rect -129 -2047 -29 -2000
rect -129 -2081 -113 -2047
rect -45 -2081 -29 -2047
rect -129 -2097 -29 -2081
rect 29 -2047 129 -2000
rect 29 -2081 45 -2047
rect 113 -2081 129 -2047
rect 29 -2097 129 -2081
<< polycont >>
rect -113 2047 -45 2081
rect 45 2047 113 2081
rect -113 -2081 -45 -2047
rect 45 -2081 113 -2047
<< locali >>
rect -289 2149 -193 2183
rect 193 2149 289 2183
rect -289 2087 -255 2149
rect 255 2087 289 2149
rect -129 2047 -113 2081
rect -45 2047 -29 2081
rect 29 2047 45 2081
rect 113 2047 129 2081
rect -175 1988 -141 2004
rect -175 -2004 -141 -1988
rect -17 1988 17 2004
rect -17 -2004 17 -1988
rect 141 1988 175 2004
rect 141 -2004 175 -1988
rect -129 -2081 -113 -2047
rect -45 -2081 -29 -2047
rect 29 -2081 45 -2047
rect 113 -2081 129 -2047
rect -289 -2149 -255 -2087
rect 255 -2149 289 -2087
rect -289 -2183 -193 -2149
rect 193 -2183 289 -2149
<< viali >>
rect -113 2047 -45 2081
rect 45 2047 113 2081
rect -175 -1988 -141 1988
rect -17 -1988 17 1988
rect 141 -1988 175 1988
rect -113 -2081 -45 -2047
rect 45 -2081 113 -2047
<< metal1 >>
rect -125 2081 -33 2087
rect -125 2047 -113 2081
rect -45 2047 -33 2081
rect -125 2041 -33 2047
rect 33 2081 125 2087
rect 33 2047 45 2081
rect 113 2047 125 2081
rect 33 2041 125 2047
rect -181 1988 -135 2000
rect -181 -1988 -175 1988
rect -141 -1988 -135 1988
rect -181 -2000 -135 -1988
rect -23 1988 23 2000
rect -23 -1988 -17 1988
rect 17 -1988 23 1988
rect -23 -2000 23 -1988
rect 135 1988 181 2000
rect 135 -1988 141 1988
rect 175 -1988 181 1988
rect 135 -2000 181 -1988
rect -125 -2047 -33 -2041
rect -125 -2081 -113 -2047
rect -45 -2081 -33 -2047
rect -125 -2087 -33 -2081
rect 33 -2047 125 -2041
rect 33 -2081 45 -2047
rect 113 -2081 125 -2047
rect 33 -2087 125 -2081
<< properties >>
string FIXED_BBOX -272 -2166 272 2166
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 20.0 l 0.5 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
